*** non-inverting amplifier ***
*global gnd
Vdd V+ 0 DC 12
Vss 0 V- DC 12
r1  0  1  1.2k
r2  1  2  43k
Vin 3 0 AC 1V
xamp1   3 1 V+ V-  2 UA741
.include UA741.cir

** Analysis setup **
.ac DEC 101 3 20.00K
.OP 
.probe
.END

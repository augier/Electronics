*** non-inverting amplifier ***
*global gnd
V1 V+ 0 DC 12
V2 0 V- DC 12
r1  0  1  1.2k
r2  1  2  9.1k
Vin 3 0 AC 1V
xamp1   3 1 V+ V-  2 UA741
.include UA741.cir

** Analysis setup **
.ac DEC 101 3 20.00K
.OP 
.probe
.END
